module TOP (
    input clk  ,
    input rst   
);
//**************************************************//
//------------------- wire define ------------------//
//**************************************************//
wire clk_lock ;
wire clk_out  ;
wire cpu_clk  ;
wire cpu_rst_n;
//**************************************************//
//--------------------- signal ---------------------//
//**************************************************//
assign cpu_clk   = clk_out & clk_lock;
assign cpu_rst_n = ~rst              ;
//**************************************************//
//--------------------- Wizard ---------------------//
//**************************************************//
CLK_Gen CLK_Gen (
    .clk_in1  ( clk      ),
    .locked   ( clk_lock ),
    .clk_out1 ( clk_out  ) 
);
//**************************************************//
//----------------------- CPU ----------------------//
//**************************************************//
RISCV RISCV (
    .clk   ( cpu_clk   ),
    .rst_n ( cpu_rst_n ) 
);

endmodule
